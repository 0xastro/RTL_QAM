--*********************************************************
---------------------------------------------------------
-- Sinsoidal Lutch 4096x12
-- Generated using Matlab
---------------------------------------------------------
-- Module: ddfs_lut_4096
-- Author: Astro
-- Project: QAM Modulation
-- Delievered to: Digital System Design
-- Supervised by: Prof. Luca Fanucci
---------------------------------------------------------
--*********************************************************

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;


ENTITY ddfs_lut_4096 is 
      port(   
            address : in std_logic_vector(11 downto 0);            -- lut address
            dds_out : out std_logic_vector(5 downto 0)             -- lut output
            );
end ddfs_lut_4096;


ARCHITECTURE bhv of ddfs_lut_4096 is
-------------------------------------------------------------------------------------
-- Internal signals & constants
-------------------------------------------------------------------------------------

TYPE int_array is ARRAY (natural range <>) of integer;            -- int_array type declaration


CONSTANT lut : int_array := (                                     -- Look up table cells/arrays
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            31,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            30,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            29,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            28,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            27,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            26,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            24,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            23,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            22,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            21,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            20,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            19,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            18,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            17,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            16,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            15,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            14,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            13,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            12,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            11,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            10,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            9,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            8,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            7,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            6,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            5,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            4,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            3,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            2,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            1,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -31,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -30,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -29,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -28,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -27,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -26,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -25,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -24,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -23,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -22,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -21,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -20,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -19,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -18,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -17,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -16,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -15,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -14,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -13,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -12,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -11,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -10,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -9,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -8,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -7,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -6,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -5,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -4,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -3,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -2,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            -1,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0);

   SIGNAL lut_address_index : integer range 0 to 4095;                              -- LUT address converted to integer to be used ad array index
      
      BEGIN
   
   lut_address_index <= to_integer(unsigned(address));                              -- Converting the lut address into an integer to be usable as array index
   
   dds_out <= std_logic_vector(to_signed(lut(lut_address_index),6));                -- Selecting the lut cell depending on the index lut_address_index

END bhv;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package arrays is
type frame is array (0 to 15) of STD_LOGIC_VECTOR;
end arrays;
